`timescale 1ns / 100ps


module pwmUnit_tb();


    /*********************************************************************************************************************************************************/
    /*                                                                                                                                                       */
    /* wire declaration                                                                                                                                      */
    /*                                                                                                                                                       */
	/*********************************************************************************************************************************************************/

	
	// input wires
    logic          clk;
	logic          reset;
	logic  [15:0]  clocksPerCycle;
	logic  [7:0]   dataIn;

	 
	// output wires
    logic          pwmOut;
	logic          readReq;

	
	/*********************************************************************************************************************************************************/
    /*                                                                                                                                                       */
    /* test module instantiation                                                                                                                             */
    /*                                                                                                                                                       */
	/*********************************************************************************************************************************************************/

    pwmUnit
	dut(
        .clk,
	    .reset,
	    .clocksPerCycle,
	    .dataIn,
	    .pwmOut,
	    .readReq
	);
	
	
	/*********************************************************************************************************************************************************/
    /*                                                                                                                                                       */
    /* testing variables                                                                                                                                     */
    /*                                                                                                                                                       */
	/*********************************************************************************************************************************************************/
	
	
	integer        seed = 125376;
	
	
	/*********************************************************************************************************************************************************/
    /*                                                                                                                                                       */
    /* test stimulus                                                                                                                                         */
    /*                                                                                                                                                       */
	/*********************************************************************************************************************************************************/
	
	
	// set initial values
	initial begin
        reset          = 1'b0;
        clocksPerCycle = 16'd8;
	    dataIn         = 8'd255;
	end
	
	
	// create clock sources
	always begin
	    #5;
	    clk = 1'b0;
	    #5;
		clk = 1'b1;
	end
	
	
	// apply test stimulus
	// synopsys translate_off
	initial begin		
		// set errors to zero
		//errorCount = 0;
		
		// set the random seed
		$urandom(seed);//x = $urandom(seed);//$srandom(seed);
		
		// reset the system
		hardwareReset();      
	
		repeat(100) begin
		    @(posedge readReq);
			@(posedge clk);
		    dataIn = $urandom();
			//@(posedge clk);
		end
		
		//$display("%d Errors", errorCount);
	    $stop;
	 end
	// synopsys translate_on

	
	/*********************************************************************************************************************************************************/
    /*                                                                                                                                                       */
    /* tasks                                                                                                                                                 */
    /*                                                                                                                                                       */
	/*********************************************************************************************************************************************************/
	
	
	task hardwareReset();
	    reset = 1'b0;
	    wait(clk !== 1'bx);
	    @(posedge clk);
	    reset = 1'b1;
	    repeat(10) @(posedge clk);
	    reset = 1'b0;
	endtask

	
endmodule

