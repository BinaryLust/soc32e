

    // uncomment this to turn on debug circuits
	//`define DEBUG

