

module vga();


// vga core clock domain 1
// contains setting registers, and font memory
// and fetches lines from memory to give to the driver

 
// vga driver clock domain 2
// receives lines from the core and drives them to the monitor


// clock domain crossing fifo


endmodule

