

package boolPkg;
	
	
    typedef enum logic {
	     T = 1'b1,
        F = 1'b0
	 }  bool;

	 
endpackage

